`ifndef soda_machine_types_sv_quard

package soda_machine_types;

	typedef enum logic [1:0] {I0=2'b00, I1=2'b01, I2=2'b10, I5=2'b11} insert_type;
	
endpackage

`define soda_machine_types_sv_quard
`endif
